// 4 BIT ADDER

module add_4_bit(a,b,sum);

    input[3:0] a,b;
    output[3:0]sum;
    
    assign sum = a + b;
    
endmodule
