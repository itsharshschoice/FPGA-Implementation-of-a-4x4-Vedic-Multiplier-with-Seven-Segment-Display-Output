// 6 BIT ADDER

module add_6_bit (a,b,sum);

    input[5:0] a,b;
    output[5:0] sum;
    
    assign sum = a + b;
    
endmodule